CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 10 5 240 9
0 66 1280 1024
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
30 D:\Program Files\CM60S\BOM.DAT
0 7
0 66 1280 1024
110100496 0
0
6 Title:
5 Name:
0
0
0
18
9 4-In AND~
219 92 285 0 5 22
0 5 2 3 4 10
0
0 0 112 90
6 74LS21
-21 -28 21 -20
4 U10A
-14 -38 14 -30
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 589832
65 0 0 0 2 1 7 0
1 U
8953 0 0
0
0
9 2-In AND~
219 194 285 0 3 22
0 9 8 11
0
0 0 112 90
6 74LS08
-21 -24 21 -16
3 U9C
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
4441 0 0
0
0
9 2-In AND~
219 161 285 0 3 22
0 9 7 12
0
0 0 112 90
6 74LS08
-21 -24 21 -16
3 U9B
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
3618 0 0
0
0
9 2-In AND~
219 127 285 0 3 22
0 9 6 13
0
0 0 112 90
6 74LS08
-21 -24 21 -16
3 U9A
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
6153 0 0
0
0
9 2-In AND~
219 402 288 0 3 22
0 6 3 19
0
0 0 112 90
6 74LS08
-21 -24 21 -16
3 U6B
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
5394 0 0
0
0
9 2-In AND~
219 352 288 0 3 22
0 2 7 20
0
0 0 112 90
6 74LS08
-21 -24 21 -16
3 U6A
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
7734 0 0
0
0
8 2-In OR~
219 372 228 0 3 22
0 20 19 21
0
0 0 112 90
6 74LS32
-21 -24 21 -16
3 U5A
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
9914 0 0
0
0
12 Hex Display~
7 372 38 0 18 19
10 2 3 4 9 0 0 0 0 0
0 1 1 1 0 1 1 1 10
0
0 0 53344 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -52 17 -44
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3747 0 0
0
0
7 Pulser~
4 28 170 0 10 12
0 23 24 22 25 0 0 5 5 4
7
0
0 0 4144 0
0
2 V1
-7 -38 7 -30
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3549 0 0
0
0
12 D Flip-Flop~
219 490 151 0 4 9
0 6 22 6 2
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 A0
-7 -58 7 -50
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
7931 0 0
0
0
12 D Flip-Flop~
219 411 151 0 4 9
0 21 22 7 3
0
0 0 5232 0
3 DFF
-10 -53 11 -45
2 U3
-7 -63 7 -55
2 A1
-6 -58 8 -50
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
9325 0 0
0
0
12 D Flip-Flop~
219 321 151 0 4 9
0 15 22 8 4
0
0 0 5232 0
3 DFF
-10 -53 11 -45
2 U2
-7 -63 7 -55
2 A2
-6 -58 8 -50
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
8903 0 0
0
0
12 D Flip-Flop~
219 240 150 0 4 9
0 14 22 5 9
0
0 0 5232 0
3 DFF
-10 -53 11 -45
2 U1
-7 -63 7 -55
2 A3
-6 -59 8 -51
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
3834 0 0
0
0
9 2-In AND~
219 281 286 0 3 22
0 4 6 18
0
0 0 112 90
6 74LS08
-21 -24 21 -16
3 U6C
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
3363 0 0
0
0
9 2-In AND~
219 315 286 0 3 22
0 4 7 17
0
0 0 112 90
6 74LS08
-21 -24 21 -16
3 U6D
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
7668 0 0
0
0
9 3-In AND~
219 246 286 0 4 22
0 8 2 3 16
0
0 0 112 90
6 74LS11
-21 -28 21 -20
3 U4A
-11 -38 10 -30
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 3 0
1 U
4718 0 0
0
0
8 3-In OR~
219 277 226 0 4 22
0 16 18 17 15
0
0 0 112 90
4 4075
-14 -24 14 -16
3 U7A
-11 -34 10 -26
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 3 5 6 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 4 0
1 U
3874 0 0
0
0
8 4-In OR~
219 137 226 0 5 22
0 10 13 12 11 14
0
0 0 112 90
4 4072
-14 -24 14 -16
3 U8A
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0
65 0 0 0 2 1 5 0
1 U
6671 0 0
0
0
42
0 2 2 0 0 4096 0 0 1 16 0 3
245 338
87 338
87 306
0 3 3 0 0 4096 0 0 1 17 0 3
254 328
96 328
96 306
0 4 4 0 0 4224 0 0 1 22 0 3
271 334
105 334
105 306
3 1 5 0 0 8320 0 13 1 0 0 6
270 132
270 171
69 171
69 310
78 310
78 306
0 2 6 0 0 4096 0 0 4 19 0 3
289 348
135 348
135 306
0 2 7 0 0 4096 0 0 3 20 0 3
324 318
169 318
169 306
0 2 8 0 0 4096 0 0 2 18 0 3
223 314
202 314
202 306
1 0 9 0 0 4096 0 2 0 0 10 2
184 306
184 324
1 0 9 0 0 0 0 3 0 0 10 2
151 306
151 324
0 1 9 0 0 12416 0 0 4 35 0 6
275 113
275 181
215 181
215 324
117 324
117 306
1 5 10 0 0 8320 0 18 1 0 0 4
127 246
127 254
91 254
91 261
4 3 11 0 0 8320 0 18 2 0 0 4
154 246
154 254
193 254
193 261
3 3 12 0 0 4224 0 18 3 0 0 3
145 246
145 261
160 261
2 3 13 0 0 4224 0 18 4 0 0 3
136 246
136 261
126 261
1 5 14 0 0 8320 0 13 18 0 0 3
216 114
140 114
140 196
0 2 2 0 0 0 0 0 16 28 0 3
342 338
245 338
245 307
0 3 3 0 0 0 0 0 16 29 0 3
411 328
254 328
254 307
3 1 8 0 0 8320 0 12 16 0 0 6
351 133
351 190
223 190
223 314
236 314
236 307
0 2 6 0 0 0 0 0 14 27 0 3
392 348
289 348
289 307
0 2 7 0 0 0 0 0 15 30 0 3
361 318
323 318
323 307
1 0 4 0 0 0 0 15 0 0 22 2
305 307
305 334
0 1 4 0 0 0 0 0 14 36 0 6
360 115
360 201
333 201
333 334
271 334
271 307
4 1 15 0 0 4224 0 17 12 0 0 3
280 196
280 115
297 115
1 4 16 0 0 8320 0 17 16 0 0 4
271 242
271 254
245 254
245 262
3 3 17 0 0 8320 0 17 15 0 0 4
289 242
289 254
314 254
314 262
2 3 18 0 0 4224 0 17 14 0 0 2
280 241
280 262
0 1 6 0 0 4224 0 0 5 34 0 4
533 133
533 348
392 348
392 309
0 1 2 0 0 4224 0 0 6 38 0 4
522 114
522 338
342 338
342 309
0 2 3 0 0 8320 0 0 5 37 0 5
450 114
451 114
451 328
410 328
410 309
3 2 7 0 0 4224 0 11 6 0 0 4
441 133
441 318
360 318
360 309
3 2 19 0 0 8320 0 5 7 0 0 4
401 264
401 259
384 259
384 244
3 1 20 0 0 8320 0 6 7 0 0 4
351 264
351 258
366 258
366 244
3 1 21 0 0 4224 0 7 11 0 0 3
375 198
375 115
387 115
3 1 6 0 0 16 0 10 10 0 0 6
520 133
533 133
533 78
460 78
460 115
466 115
4 4 9 0 0 0 0 8 13 0 0 5
363 62
363 69
275 69
275 114
264 114
3 4 4 0 0 0 0 8 12 0 0 5
369 62
369 78
360 78
360 115
345 115
2 4 3 0 0 0 0 8 11 0 0 5
375 62
375 78
450 78
450 115
435 115
1 4 2 0 0 0 0 8 10 0 0 5
381 62
381 68
522 68
522 115
514 115
2 0 22 0 0 8192 0 13 0 0 42 3
216 132
210 132
210 161
2 0 22 0 0 0 0 12 0 0 42 3
297 133
290 133
290 161
2 0 22 0 0 0 0 11 0 0 42 3
387 133
382 133
382 161
3 2 22 0 0 4224 0 9 10 0 0 4
52 161
462 161
462 133
466 133
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
